�� sr Repositories.TestingTableRepo      � L testingTableListt Ljava/util/List;xpsr java.util.ArrayListx����a� I sizexp   w   sr domains.TestingTable      � J 	studentIdJ 	variantIdxp              sq ~               sq ~               sq ~               sq ~               x