�� sr Repositories.VariantsRepo      � J elementsCountJ 
idSequenceL variantsListt Ljava/util/List;xp              sr java.util.ArrayListx����a� I sizexp   w   sr domains.Variant      � J idL 
pathToFilet Ljava/lang/String;xp       t var1sq ~        t var7sq ~        t var2sq ~        t var3sq ~        t var4sq ~        t var5sq ~        t var6x