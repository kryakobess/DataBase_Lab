�� sr Repositories.StudentsRepo      � J elementsCountJ 
idSequenceL studentsListt Ljava/util/List;xp       ^       ^sr java.util.ArrayListx����a� I sizexp   ^w   ^sr domains.Student      � J idL namet Ljava/lang/String;L 
patronymicq ~ L surnameq ~ xp       t Максимt Александровичt 
Агеевsq ~        t Андрейt Николаевичt Акимовsq ~        t Максимt Сергеевичt Анохинsq ~        t Юрийt Валерьевичt Антиповsq ~        t Дмитрийt Алексеевичt Антоновsq ~        t Богданt Михайловичt Артемьевsq ~        t Кириллt Ивановичt 
Бабинsq ~        t Матвейt 
Ильичt Барышевsq ~        	t Андрейt Сергеевичt Безуховsq ~        
t Светланаt Евгеньевнаt Болотинаsq ~        t Елизаветаt Юрьевнаt Борисоваsq ~        t Дастанt Маратовичt Буларкиевsq ~        t 
Дарьяt Григорьевнаt Вавиловаsq ~        t Олегt Александровичt 
Вагинsq ~        t Анастасияt Георгиевнаt Вайнерsq ~        t Данилаt Валерьевичt Веряскинsq ~        t Владиславt Сергеевичt Волковsq ~        t Филиппt Олеговичt Волковsq ~        t Ильяt Сергеевичt Володинsq ~        t Надеждаt Артемовнаt Воропаеваsq ~        t Сергейt Николаевичt Горячевsq ~        t Николайt Алексеевичt Грызловsq ~        t Русланt -t Даминовsq ~        t Егорt Васильевичt Дементьевsq ~        t Ильяt Михайловичt Доманскийsq ~        t Максимt Александровичt Дударевsq ~        t Елизаветаt Андреевнаt Захароваsq ~        t Анатолийt Максимовичt Иванашкоsq ~        t 
Данилt Вадимовичt Калининsq ~        t 
Игорьt Александровичt Камышенковsq ~        t 
Элинаt Камоевнаt Карапетянsq ~         t 
Вадимt Александровичt Карповsq ~        !t Анастасияt -t Катауроваsq ~        "t Екатеринаt -t Кенегесоваsq ~        #t Ильяt Сергеевичt Кобызевsq ~        $t 
Борисt Алексеевичt 
Козинsq ~        %t Иванt Федоровичt Коломинскийsq ~        &t Юлияt Андреевнаt Комароваsq ~        't Зояt Константиновнаt Кораблеваsq ~        (t Ильяt Андреевичt Кравченкоsq ~        )t Серафимt Павловичt Кравчукsq ~        *t Ильяt Михайловичt Крамникsq ~        +t Иванt Владимировичt Курихинsq ~        ,t Никитаt Александровичt Курицынsq ~        -t Владиславt Сергеевичt Курылевsq ~        .t Дмитрийt Николаевичt Кутузовsq ~        /t 
Ольгаt Александровнаt Лакееваsq ~        0t 
Игорьt -t Мамонтовsq ~        1t 
Павелt Александровичt Медведевsq ~        2t Маринаt Васильевнаt Мельникsq ~        3t Максимt Дмитриевичt Молчановsq ~        4t 
Артёмt Вадимовичt Муштуковsq ~        5t 
Аленаt Алексеевнаt Нишнючкинаsq ~        6t Ильяt Павловичt Носковsq ~        7t 
Алинаt Андреевнаt Обрезковаsq ~        8t Евгенийt Данииловичt Парфененковsq ~        9t 
Антонt -t Пестриковsq ~        :t Дмитрийt Андреевичt Петровsq ~        ;t Андрейt Владимировичt Помошниковsq ~        <t Станиславt Игоревичt Романовsq ~        =t Андрейt Дмитриевичt 
Рябовsq ~        >t Максимt Александровичt Саляевsq ~        ?t Максимt Вячеславовичt Селезневsq ~        @t Никитаt Сергеевичt Семеновsq ~        At 
Олесяt Николаевнаt Сергееваsq ~        Bt 
Марияt Игоревнаt Симоноваsq ~        Ct 
Марияt Дмитриевнаt Слепневаsq ~        Dt 
Алинаt Денисовнаt Сологубsq ~        Et Даниилt Дмитриевичt Солынинsq ~        Ft Русланt Наримановичt Сорокинsq ~        Gt Всеволодt 
Ильичt Сорокинsq ~        Ht Иванt Александровичt Стасевичsq ~        It Максимt Олеговичt Столетовsq ~        Jt Петрt Викторовичt Стрельниковsq ~        Kt Русланt Аликовичt Султановsq ~        Lt Василийt Андреевичt Сунцовsq ~        Mt Алексейt Олеговичt Талановsq ~        Nt Пётрt Вячеславовичt Тюхменевsq ~        Ot Отабекt Айбековичt Уразмахатовsq ~        Pt Екатеринаt Владимировнаt Уржумцеваsq ~        Qt Эдемt Икромовичt Хадиевsq ~        Rt Натальяt Васильевнаt Христолюбоваsq ~        St Георгийt Максимовичt Чайкинsq ~        Tt Алексейt Владимировичt Черепановsq ~        Ut Михаилt Алексеевичt Чернышевскийsq ~        Vt 
Антонt Альбертовичt Шадринsq ~        Wt Андрейt Сергеевичt 
Шаровsq ~        Xt Юлияt Юрьевнаt Шаталинаsq ~        Yt 
Романt Андреевичt Шемановскийsq ~        Zt 
Данилt Сергеевичt Шероновsq ~        [t 
Эрикаt Лунаt 
Шиминsq ~        \t Юрийt Игоревичt 
Шоринsq ~        ]t Данилаt Андреевичt Шуваевsq ~        ^t Владиславt Юрьевичt Щегловx