�� sr Repositories.StudentsRepo      � J elementsCountJ 
idSequenceL studentsListt Ljava/util/List;xp              sr java.util.ArrayListx����a� I sizexp   w   sr domains.Student      � J idL namet Ljava/lang/String;L 
patronymicq ~ L surnameq ~ xp       t Nikitat Alext Kuritsynsq ~        t Bubat  t Bibasq ~        t Kuritaq ~ 	t 
Nikititsynsq ~        t hehet bebet huhusq ~        q ~ q ~ t Bebax